library IEEE;
use 	IEEE.STD_LOGIC_1164.ALL;
use 	IEEE.STD_LOGIC_ARITH.ALL;
use 	IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Sumador1bit is
	port (A : in STD_LOGIC;
			B : in STD_LOGIC;
			C_in : STD_LOGIC;
			Suma : out STD_LOGIC;
			Acarreo : out STD_LOGIC;
end Sumador1bit;

architecture behavior of Sumador1bit is
end behavior;

